
module keyBounce(
	input logic [3:0] decoded key
);


endmodule
